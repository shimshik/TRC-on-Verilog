module driver7seg (
input[3:0] bin,
output[6*7-1:0] hex
);
reg [6*7-1:0] rhex;
always@*
case(bin)
4'b0000: rhex=42'b1111111_1111111_1111111_0000010_1000000_0001100; // GoToWork
4'b0001: rhex=42'b1111111_1111111_1111111_1111111_0010010_0001100; // StopWork
4'b0010: rhex=42'b1111111_1111111_1111111_1111111_0000010_0010010; // GoToSt
4'b0011: rhex=42'b1111111_1111111_1111111_0001000_1111011_0000111; // Wait
4'b0100: rhex=42'b1111111_1111111_1111111_1111111_0100001_1000000; // DrsIsOpen
4'b0101: rhex=42'b1111111_1111111_1111111_0100001_1000110_1000000; // DrsCntOpen
4'b0110: rhex=42'b1111111_1111111_1111111_1111111_0100001_1000110; // DrsIsClose
4'b0111: rhex=42'b1111111_1111111_1111111_0100001_1000110_1000110; // DrsCntClose
4'b1000: rhex=42'b1111111_0000110_0101111_0101111_1000000_0101111; // SmthWrong



endcase
assign hex=rhex;
endmodule
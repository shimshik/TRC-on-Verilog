// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus II Version 15.0.0 Build 145 04/22/2015 SJ Web Edition
// Created on Wed Dec 18 18:00:33 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module moore (
    reset,clock,ctrl,
    evnt[3:0]);

    input reset;
    input clock;
    input ctrl;
    tri0 reset;
    tri0 ctrl;
    output [3:0] evnt;
    reg [3:0] evnt;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter START=0,A=1,B=2,C=3,D=4;

    always @(posedge clock or negedge reset)
    begin
        if (~reset) begin
            fstate <= START;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or ctrl)
    begin
        evnt <= 4'b0000;
        case (fstate)
            START: begin
                if (ctrl)
                    reg_fstate <= C;
                else if (~(ctrl))
                    reg_fstate <= A;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= START;

                evnt <= 4'b0000;
            end
            A: begin
                if (ctrl)
                    reg_fstate <= A;
                else if (~(ctrl))
                    reg_fstate <= B;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= A;

                evnt <= 4'b0001;
            end
            B: begin
                if (ctrl)
                    reg_fstate <= B;
                else if (~(ctrl))
                    reg_fstate <= C;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= B;

                evnt <= 4'b0010;
            end
            C: begin
                reg_fstate <= D;

                evnt <= 4'b0011;
            end
            D: begin
                if (ctrl)
                    reg_fstate <= C;
                else if (~(ctrl))
                    reg_fstate <= D;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= D;

                evnt <= 4'b0100;
            end
            default: begin
                evnt <= 4'bxxxx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // moore
